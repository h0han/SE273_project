----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2020/11/27 23:56:15
-- Design Name: 
-- Module Name: SEVENBIT_ADDER - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SEVENBIT_ADDER is
    Port ( A : in STD_LOGIC_VECTOR (6 downto 0);
           B : in STD_LOGIC_VECTOR (6 downto 0);
           C : out STD_LOGIC_VECTOR (6 downto 0));
end SEVENBIT_ADDER;

architecture Behavioral of SEVENBIT_ADDER is

begin


end Behavioral;
